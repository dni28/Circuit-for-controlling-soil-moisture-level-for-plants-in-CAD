** Profile: "SCHEMATIC1-DC_Sweep2"  [ C:\Users\salaj\Desktop\Proiect_CAD\Project_CAD-PSpiceFiles\SCHEMATIC1\DC_Sweep2.sim ] 

** Creating circuit file "DC_Sweep2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Cadence_Orcad\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM rvar 600k 60k -1k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
